//non-parameterized class extended from non-parameterized class
