`include "parameterized_memory.v"
`include "mem_intf.sv"
`include "mem_common.sv"
`include "mem_tx.sv"
//`include "mem_bfm.sv"
`include "mem_bfm_cb_mp.sv"
`include "mem_gen.sv"
`include "mem_mon.sv"
`include "mem_cov.sv"
`include "mem_agent.sv"
`include "mem_env.sv"
`include "tb_top.sv"

