class mem_env;
mem_agent agent = new();
	
task run();
	agent.run();
endtask
	
endclass