class eth_pkt_common;
	static mailbox gen2bfm_mb = new(); //common mailbox between generator and driver/bfm.
	static string test_case_name;
	static integer no_of_packets = 20;
endclass