//wild card operators - some positions in the vector, we don't want to check, it doesn't matter whether  that bit is 1 or 0,
//that specific position check will be ignored.
// (a==?b) --> if b has any x or z, those positions will not be compared. 
//-But if 'a' has x or z --> output of comaprison will be 'x'.

module tb;



endmodule 
