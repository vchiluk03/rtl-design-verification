library verilog;
use verilog.vl_types.all;
entity tb is
    generic(
        WIDTH_TB        : integer := 15
    );
end tb;
