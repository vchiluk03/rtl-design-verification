library verilog;
use verilog.vl_types.all;
entity tb is
    generic(
        NUM             : integer := 9
    );
end tb;
